//**********************************************
//**********    gatelevel module   *************

    // ----------------------   
    //  FILL YOUR CODE HERE
    // ----------------------
